`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: NUS
// Engineer: Shahzor Ahmad, Rajesh C Panicker
// 
// Create Date: 27.09.2016 10:59:44
// Design Name: 
// Module Name: MCycle
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
/* 
----------------------------------------------------------------------------------
--	(c) Shahzor Ahmad, Rajesh C Panicker
--	License terms :
--	You are free to use this code as long as you
--		(i) DO NOT post it on any public repository;
--		(ii) use it only for educational purposes;
--		(iii) accept the responsibility to ensure that your implementation does not violate any intellectual property of ARM Holdings or other entities.
--		(iv) accept that the program is provided "as is" without warranty of any kind or assurance regarding its suitability for any particular purpose;
--		(v) send an email to rajesh.panicker@ieee.org briefly mentioning its use (except when used for the course CG3207 at the National University of Singapore);
--		(vi) retain this notice in this file or any files derived from this.
----------------------------------------------------------------------------------
*/

module MCycle

    #(parameter width = 4) // Keep this at 4 to verify your algorithms with 4 bit numbers (easier). When using MCycle as a component in ARM, generic map it to 32.
    (
        input CLK,
        input RESET, // Connect this to the reset of the ARM processor.
        input Start, // Multi-cycle Enable. The control unit should assert this when an instruction with a multi-cycle operation is detected.
        input [1:0] MCycleOp, // Multi-cycle Operation. "00" for signed multiplication, "01" for unsigned multiplication, "10" for signed division, "11" for unsigned division. Generated by Control unit
        input [width-1:0] Operand1, // Multiplicand / Dividend
        input [width-1:0] Operand2, // Multiplier / Divisor
        output reg [width-1:0] Result1, // LSW of Product / Quotient
        output reg [width-1:0] Result2, // MSW of Product / Remainder
        output reg Busy // Set immediately when Start is set. Cleared when the Results become ready. This bit can be used to stall the processor while multi-cycle operations are on.
    );
    
// use the Busy signal to reset WE_PC to 0 in ARM.v (aka "freeze" PC). The two signals are complements of each other
// since the IDLE_PROCESS is combinational, instantaneously asserts Busy once Start is asserted
  
    parameter IDLE = 1'b0 ;  // will cause a warning which is ok to ignore - [Synth 8-2507] parameter declaration becomes local in MCycle with formal parameter declaration list...

    parameter COMPUTING = 1'b1 ; // this line will also cause the above warning
    reg state = IDLE ;
    reg n_state = IDLE ;
   
    reg [7:0] count = 0 ; // assuming no computation takes more than 256 cycles.
    
    reg done;
    
    // Multiplication related registers
    reg [2*width-1:0] temp_sum = 0 ;        // accumulator for multiplication
    reg [2*width-1:0] temp_sum_after_op;  
    reg [2*width-1:0] shifted_op1_mul = 0 ; // multiplicand
    reg [width-1:0] shifted_op2_mul = 0 ; // multiplier   
    reg carry = 0 ;
    reg [1:0] qn = 0;

    // Division related registers
    reg [2*width:0] op2_abs; // Absolute value of Divisor
    reg quotient_sign;
    reg remainder_sign;
    reg [width-1:0] quotient_abs;
    reg [2*width:0] remainder_abs;
    reg [2*width:0] temp_remainder;
    
    always@( state, done, Start, RESET ) begin : IDLE_PROCESS  
		// Note : This block uses non-blocking assignments to get around an unpredictable Verilog simulation behaviour.
        // default outputs
        Busy <= 1'b0 ;
        n_state <= IDLE ;
        
        // reset
        if(~RESET)
            case(state)
                IDLE: begin
                    if(Start) begin // note: a mealy machine, since output depends on current state (IDLE) & input (Start)
                        n_state <= COMPUTING ;
                        Busy <= 1'b1 ;
                    end
                end
                COMPUTING: begin
                    if(~done) begin
                        n_state <= COMPUTING ;
                        Busy <= 1'b1 ;
                    end
                end        
            endcase    
    end


    always@( posedge CLK ) begin : STATE_UPDATE_PROCESS // state updating
        state <= n_state ;    
    end

    
    always@( posedge CLK ) begin : COMPUTING_PROCESS // process which does the actual computation
        // n_state == COMPUTING and state == IDLE implies we are just transitioning into COMPUTING
        if( RESET | (n_state == COMPUTING & state == IDLE) ) begin // 2nd condition is true during the very 1st clock cycle of the multiplication
            count <= 0;
            done <= 1'b0 ;

            // Multiplication initialisation
            temp_sum <= 0 ;
            
            if (MCycleOp == 2'b00) begin // Signed Multiplication
                shifted_op1_mul <= Operand1[width-1] ? {{(width+1){1'b1}}, Operand1} : {{(width+1){1'b0}}, Operand1}; // sign/zero extend the operands
                shifted_op2_mul <= Operand2;
                carry <= 1'b0;
            end else if (MCycleOp == 2'b01) begin // Unsigned Multiplication
                shifted_op1_mul <= {{(width){1'b0}}, Operand1};
                shifted_op2_mul <= Operand2;
            end

            // Division initialisation
            else if (MCycleOp == 2'b10) begin // Signed Division
                remainder_abs <= Operand1[width-1] ? {{(width+1){1'b0}}, ~Operand1 + 1'b1} : {{(width+1){1'b0}}, Operand1};
                op2_abs <= Operand2[width-1] ? {1'b0, (~Operand2 + 1'b1), {width{1'b0}}} : {1'b0, Operand2, {{width{1'b0}}}}; // absolute value of Divisor
                quotient_sign <= Operand1[width-1] ^ Operand2[width-1]; // sign of Quotient
                remainder_sign <= Operand1[width-1]; // sign of Remainder = sign of Dividend
                quotient_abs <= 1'b0;
            end else begin // Unsigned Division
                remainder_abs <= {{(width+1){1'b0}}, Operand1};
                op2_abs <= {1'b0, Operand2, {{width{1'b0}}}};
                quotient_sign <= 1'b0;
                remainder_sign <= 1'b0;
                quotient_abs <= 1'b0;
            end

            Result1 <= 0 ;
            Result2 <= 0 ;
        end 

        else if (state == COMPUTING) begin
            count <= count + 1;
            done <= 1'b0 ;

            if (MCycleOp == 2'b01) begin // Unsigned multiplication 
                if(shifted_op2_mul[0]) // add only if LSB of multiplier is 1
                temp_sum = temp_sum + shifted_op1_mul ; // partial product for multiplication
                
                shifted_op2_mul = {1'b0, shifted_op2_mul[width-1 : 1]} ;
                shifted_op1_mul = {shifted_op1_mul[2*width-2 : 0], 1'b0} ; 

                if (count == width-1)
                    done <= 1'b1 ; 

                Result2 <= temp_sum[2*width-1 : width] ;
                Result1 <= temp_sum[width-1 : 0] ; 
            end else if (MCycleOp == 2'b00) begin
               // Booth's algorithm for signed multiplication
               qn = {shifted_op2_mul[0], carry};
               
               case(qn)
                   2'b01:  temp_sum_after_op = temp_sum + shifted_op1_mul;      // A = A + M
                   2'b10:  temp_sum_after_op = temp_sum - shifted_op1_mul;      // A = A - M
                   default: temp_sum_after_op = temp_sum;                       // No operation
               endcase

               carry <= shifted_op2_mul[0];
               shifted_op2_mul <= {temp_sum_after_op[0], shifted_op2_mul[width-1:1]}; 
               temp_sum <= {temp_sum_after_op[2*width-1], temp_sum_after_op[2*width-1:1]}; 

               if (count == width) 
                   done <= 1'b1 ;           

               Result2 <= temp_sum[width-1:0] ;      
               Result1 <= shifted_op2_mul;
            end else begin // Divide
                temp_remainder = remainder_abs + ~op2_abs + 1'b1;
                if (temp_remainder[2*width]) begin // remainder < divisor
                    quotient_abs <= {quotient_abs[width-2:0], 1'b0};
                end else begin
                    remainder_abs <= temp_remainder;
                    quotient_abs <= {quotient_abs[width-2:0], 1'b1};
                end
                
                op2_abs <= {1'b0, op2_abs[2*width:1]};
                
                if (count == width + 1) begin
                    done <= 1'b1;
                end
                
                Result1 <= quotient_sign ? ~quotient_abs + 1'b1 : quotient_abs;
                Result2 <= remainder_sign ? ~remainder_abs[width-1:0] + 1'b1 : remainder_abs[width-1:0];
            end
        end
    end
endmodule